LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

ENTITY function_81 IS
    PORT (
        --missing
    );
END function_81;

ARCHITECTURE rtl OF function_81 IS

    COMPONENT mux81 IS
        PORT (
            i1_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            i2_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            i3_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            i4_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            i5_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            i6_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            i7_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            i8_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            sel_81 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            y_81 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
    END COMPONENT mux81;

BEGIN
    --missing
END rtl;