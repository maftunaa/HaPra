library ieee;
use ieee.std_logic_1164.all;

entity ms_ff is
    port (
      d, clk: in std_logic;
      Q, not_Q : out std_logic
    );
  end ms_ff;

architecture behavioral of ms_ff is

--missing

--missing

begin

--missing

end behavioral ;