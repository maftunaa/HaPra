library ieee;
use ieee.std_logic_1164.all;

entity D_Latch is
    port(
        D, clk : in std_logic;
        Q, not_Q : out std_logic
    );
end D_Latch;

architecture Behavioral of D_Latch is
    
--missing

begin

--missing

end Behavioral;