library ieee;
use ieee.std_logic_1164.all;

entity ms_ff_tb is
end ms_ff_tb;

architecture testbench of ms_ff_tb is

--missing

begin
   
--missing
   
end testbench;