library ieee;
use ieee.std_logic_1164.all;

entity ff_reset_tb is
end ff_reset_tb;

architecture testbench of ff_reset_tb is

--missing

begin
   
--missing
   
end testbench;