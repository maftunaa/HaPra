library ieee;
use ieee.std_logic_1164.all;

entity ff_reset is
    port (
      d, clk, reset: in std_logic;
      Q, not_Q : out std_logic
    );
  end ff_reset;

architecture behavioral of ff_reset is

--missing

--missing

begin

--missing

end behavioral ;